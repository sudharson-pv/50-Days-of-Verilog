module decoder3_8(input [2:0] a, output [7:0] y);
    assign y = 8'b00000001 << a;
endmodule




